VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1429.100 2924.800 1430.300 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2228.650 3517.600 2229.210 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.810 3517.600 1905.370 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.970 3517.600 1581.530 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.290 3517.600 933.850 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.450 3517.600 610.010 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.610 3517.600 286.170 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3471.140 2.400 3472.340 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3212.740 2.400 3213.940 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2954.340 2.400 2955.540 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1692.940 2924.800 1694.140 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2695.940 2.400 2697.140 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2437.540 2.400 2438.740 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2179.140 2.400 2180.340 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1920.740 2.400 1921.940 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1662.340 2.400 1663.540 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1403.940 2.400 1405.140 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1145.540 2.400 1146.740 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 887.140 2.400 888.340 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 628.740 2.400 629.940 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1956.780 2924.800 1957.980 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2220.620 2924.800 2221.820 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2484.460 2924.800 2485.660 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2748.300 2924.800 2749.500 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3012.140 2924.800 3013.340 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3275.980 2924.800 3277.180 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2876.330 3517.600 2876.890 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2552.490 3517.600 2553.050 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 43.940 2924.800 45.140 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2286.580 2924.800 2287.780 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2550.420 2924.800 2551.620 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2814.260 2924.800 2815.460 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.100 2924.800 3079.300 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3341.940 2924.800 3343.140 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2795.370 3517.600 2795.930 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2471.530 3517.600 2472.090 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2147.690 3517.600 2148.250 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1823.850 3517.600 1824.410 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.010 3517.600 1500.570 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 241.820 2924.800 243.020 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.170 3517.600 1176.730 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.330 3517.600 852.890 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.490 3517.600 529.050 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.650 3517.600 205.210 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3406.540 2.400 3407.740 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3148.140 2.400 3149.340 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2889.740 2.400 2890.940 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2631.340 2.400 2632.540 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2372.940 2.400 2374.140 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2114.540 2.400 2115.740 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 439.700 2924.800 440.900 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1856.140 2.400 1857.340 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1597.740 2.400 1598.940 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1339.340 2.400 1340.540 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1080.940 2.400 1082.140 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 822.540 2.400 823.740 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 564.140 2.400 565.340 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 370.340 2.400 371.540 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 176.540 2.400 177.740 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 637.580 2924.800 638.780 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 835.460 2924.800 836.660 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1033.340 2924.800 1034.540 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1231.220 2924.800 1232.420 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1495.060 2924.800 1496.260 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1758.900 2924.800 1760.100 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2022.740 2924.800 2023.940 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 175.860 2924.800 177.060 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2418.500 2924.800 2419.700 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2682.340 2924.800 2683.540 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2946.180 2924.800 2947.380 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3210.020 2924.800 3211.220 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3473.860 2924.800 3475.060 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2633.450 3517.600 2634.010 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2309.610 3517.600 2310.170 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1985.770 3517.600 1986.330 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.930 3517.600 1662.490 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 373.740 2924.800 374.940 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.250 3517.600 1014.810 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.410 3517.600 690.970 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.570 3517.600 367.130 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.730 3517.600 43.290 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3277.340 2.400 3278.540 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3018.940 2.400 3020.140 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2760.540 2.400 2761.740 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2502.140 2.400 2503.340 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2243.740 2.400 2244.940 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1985.340 2.400 1986.540 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 571.620 2924.800 572.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1726.940 2.400 1728.140 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1468.540 2.400 1469.740 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1210.140 2.400 1211.340 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 951.740 2.400 952.940 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 693.340 2.400 694.540 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 434.940 2.400 436.140 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 241.140 2.400 242.340 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 47.340 2.400 48.540 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 769.500 2924.800 770.700 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1165.260 2924.800 1166.460 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1363.140 2924.800 1364.340 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1626.980 2924.800 1628.180 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1890.820 2924.800 1892.020 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2154.660 2924.800 2155.860 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 109.900 2924.800 111.100 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2352.540 2924.800 2353.740 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2616.380 2924.800 2617.580 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2880.220 2924.800 2881.420 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3144.060 2924.800 3145.260 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3407.900 2924.800 3409.100 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2714.410 3517.600 2714.970 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.570 3517.600 2391.130 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2066.730 3517.600 2067.290 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.890 3517.600 1743.450 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 307.780 2924.800 308.980 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.210 3517.600 1095.770 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.370 3517.600 771.930 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.530 3517.600 448.090 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.690 3517.600 124.250 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3341.940 2.400 3343.140 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3083.540 2.400 3084.740 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2825.140 2.400 2826.340 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2566.740 2.400 2567.940 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2308.340 2.400 2309.540 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2049.940 2.400 2051.140 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 505.660 2924.800 506.860 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1791.540 2.400 1792.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1533.140 2.400 1534.340 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1274.740 2.400 1275.940 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1016.340 2.400 1017.540 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 757.940 2.400 759.140 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 499.540 2.400 500.740 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 305.740 2.400 306.940 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 111.940 2.400 113.140 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 703.540 2924.800 704.740 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 901.420 2924.800 902.620 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1099.300 2924.800 1100.500 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1297.180 2924.800 1298.380 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1561.020 2924.800 1562.220 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1824.860 2924.800 1826.060 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2088.700 2924.800 2089.900 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.970 -4.800 684.530 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2339.970 -4.800 2340.530 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2356.530 -4.800 2357.090 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2373.090 -4.800 2373.650 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2389.650 -4.800 2390.210 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2406.210 -4.800 2406.770 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2439.330 -4.800 2439.890 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2455.890 -4.800 2456.450 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2472.450 -4.800 2473.010 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2489.010 -4.800 2489.570 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.570 -4.800 850.130 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2505.570 -4.800 2506.130 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2522.130 -4.800 2522.690 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.690 -4.800 2539.250 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2555.250 -4.800 2555.810 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2588.370 -4.800 2588.930 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2604.930 -4.800 2605.490 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.490 -4.800 2622.050 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.050 -4.800 2638.610 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2654.610 -4.800 2655.170 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.130 -4.800 866.690 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2671.170 -4.800 2671.730 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2687.730 -4.800 2688.290 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2704.290 -4.800 2704.850 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2720.850 -4.800 2721.410 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2737.410 -4.800 2737.970 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2753.970 -4.800 2754.530 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2770.530 -4.800 2771.090 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2787.090 -4.800 2787.650 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.250 -4.800 899.810 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.810 -4.800 916.370 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 -4.800 932.930 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.930 -4.800 949.490 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.490 -4.800 966.050 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.050 -4.800 982.610 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.610 -4.800 999.170 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.530 -4.800 701.090 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.170 -4.800 1015.730 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.730 -4.800 1032.290 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.290 -4.800 1048.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.850 -4.800 1065.410 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.410 -4.800 1081.970 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.970 -4.800 1098.530 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.090 -4.800 1131.650 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.650 -4.800 1148.210 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.210 -4.800 1164.770 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.090 -4.800 717.650 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.770 -4.800 1181.330 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.330 -4.800 1197.890 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1213.890 -4.800 1214.450 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.450 -4.800 1231.010 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.010 -4.800 1247.570 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.570 -4.800 1264.130 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.130 -4.800 1280.690 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1296.690 -4.800 1297.250 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.250 -4.800 1313.810 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.810 -4.800 1330.370 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.650 -4.800 734.210 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.930 -4.800 1363.490 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.490 -4.800 1380.050 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.050 -4.800 1396.610 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1412.610 -4.800 1413.170 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.170 -4.800 1429.730 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.730 -4.800 1446.290 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.290 -4.800 1462.850 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.850 -4.800 1479.410 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.210 -4.800 750.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1511.970 -4.800 1512.530 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1528.530 -4.800 1529.090 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.650 -4.800 1562.210 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1578.210 -4.800 1578.770 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1594.770 -4.800 1595.330 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.330 -4.800 1611.890 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1644.450 -4.800 1645.010 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.010 -4.800 1661.570 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.770 -4.800 767.330 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1677.570 -4.800 1678.130 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1694.130 -4.800 1694.690 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.810 -4.800 1744.370 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.370 -4.800 1760.930 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.930 -4.800 1777.490 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.050 -4.800 1810.610 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1826.610 -4.800 1827.170 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.330 -4.800 783.890 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1843.170 -4.800 1843.730 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1859.730 -4.800 1860.290 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1892.850 -4.800 1893.410 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1909.410 -4.800 1909.970 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1925.970 -4.800 1926.530 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1942.530 -4.800 1943.090 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1975.650 -4.800 1976.210 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1992.210 -4.800 1992.770 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.890 -4.800 800.450 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2008.770 -4.800 2009.330 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2025.330 -4.800 2025.890 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2058.450 -4.800 2059.010 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2075.010 -4.800 2075.570 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2091.570 -4.800 2092.130 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2108.130 -4.800 2108.690 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2141.250 -4.800 2141.810 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2157.810 -4.800 2158.370 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.450 -4.800 817.010 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2174.370 -4.800 2174.930 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.050 -4.800 2224.610 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2240.610 -4.800 2241.170 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2257.170 -4.800 2257.730 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2273.730 -4.800 2274.290 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2306.850 -4.800 2307.410 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2323.410 -4.800 2323.970 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.010 -4.800 833.570 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.490 -4.800 690.050 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2362.050 -4.800 2362.610 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2395.170 -4.800 2395.730 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2411.730 -4.800 2412.290 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2428.290 -4.800 2428.850 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2444.850 -4.800 2445.410 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2477.970 -4.800 2478.530 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.090 -4.800 855.650 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2511.090 -4.800 2511.650 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2527.650 -4.800 2528.210 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2560.770 -4.800 2561.330 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2577.330 -4.800 2577.890 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2593.890 -4.800 2594.450 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2610.450 -4.800 2611.010 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2643.570 -4.800 2644.130 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2660.130 -4.800 2660.690 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.650 -4.800 872.210 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2676.690 -4.800 2677.250 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2693.250 -4.800 2693.810 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2742.930 -4.800 2743.490 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2759.490 -4.800 2760.050 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2776.050 -4.800 2776.610 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.210 -4.800 888.770 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.770 -4.800 905.330 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.330 -4.800 921.890 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.890 -4.800 938.450 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.450 -4.800 955.010 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.010 -4.800 971.570 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.570 -4.800 988.130 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.130 -4.800 1004.690 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.050 -4.800 706.610 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.690 -4.800 1021.250 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.810 -4.800 1054.370 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.370 -4.800 1070.930 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.930 -4.800 1087.490 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1103.490 -4.800 1104.050 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.050 -4.800 1120.610 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.610 -4.800 1137.170 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1153.170 -4.800 1153.730 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.730 -4.800 1170.290 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.610 -4.800 723.170 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.290 -4.800 1186.850 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.850 -4.800 1203.410 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1219.410 -4.800 1219.970 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1235.970 -4.800 1236.530 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.530 -4.800 1253.090 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.650 -4.800 1286.210 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.210 -4.800 1302.770 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.770 -4.800 1319.330 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.330 -4.800 1335.890 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.170 -4.800 739.730 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1351.890 -4.800 1352.450 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.450 -4.800 1369.010 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.010 -4.800 1385.570 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.570 -4.800 1402.130 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1434.690 -4.800 1435.250 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.250 -4.800 1451.810 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.810 -4.800 1468.370 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.370 -4.800 1484.930 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.930 -4.800 1501.490 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.730 -4.800 756.290 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.490 -4.800 1518.050 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.050 -4.800 1534.610 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.610 -4.800 1551.170 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1567.170 -4.800 1567.730 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.730 -4.800 1584.290 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.290 -4.800 1600.850 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.850 -4.800 1617.410 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.410 -4.800 1633.970 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1666.530 -4.800 1667.090 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.290 -4.800 772.850 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.090 -4.800 1683.650 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.650 -4.800 1700.210 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.210 -4.800 1716.770 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.770 -4.800 1733.330 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.330 -4.800 1749.890 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1765.890 -4.800 1766.450 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1782.450 -4.800 1783.010 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.010 -4.800 1799.570 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1815.570 -4.800 1816.130 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1832.130 -4.800 1832.690 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.850 -4.800 789.410 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1848.690 -4.800 1849.250 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1865.250 -4.800 1865.810 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1898.370 -4.800 1898.930 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1914.930 -4.800 1915.490 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1931.490 -4.800 1932.050 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1948.050 -4.800 1948.610 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1964.610 -4.800 1965.170 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1981.170 -4.800 1981.730 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1997.730 -4.800 1998.290 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2014.290 -4.800 2014.850 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.850 -4.800 2031.410 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.410 -4.800 2047.970 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2063.970 -4.800 2064.530 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.530 -4.800 2081.090 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2097.090 -4.800 2097.650 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.210 -4.800 2130.770 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2146.770 -4.800 2147.330 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2163.330 -4.800 2163.890 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.970 -4.800 822.530 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2179.890 -4.800 2180.450 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2196.450 -4.800 2197.010 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2229.570 -4.800 2230.130 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2246.130 -4.800 2246.690 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2262.690 -4.800 2263.250 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2279.250 -4.800 2279.810 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2312.370 -4.800 2312.930 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.930 -4.800 2329.490 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.530 -4.800 839.090 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.010 -4.800 695.570 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2351.010 -4.800 2351.570 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.570 -4.800 2368.130 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.130 -4.800 2384.690 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2400.690 -4.800 2401.250 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2433.810 -4.800 2434.370 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2450.370 -4.800 2450.930 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2466.930 -4.800 2467.490 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2483.490 -4.800 2484.050 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2500.050 -4.800 2500.610 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.610 -4.800 861.170 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2516.610 -4.800 2517.170 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2533.170 -4.800 2533.730 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2549.730 -4.800 2550.290 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2566.290 -4.800 2566.850 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2582.850 -4.800 2583.410 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2599.410 -4.800 2599.970 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2615.970 -4.800 2616.530 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.530 -4.800 2633.090 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2665.650 -4.800 2666.210 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2682.210 -4.800 2682.770 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2698.770 -4.800 2699.330 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2715.330 -4.800 2715.890 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2731.890 -4.800 2732.450 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2748.450 -4.800 2749.010 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2765.010 -4.800 2765.570 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2781.570 -4.800 2782.130 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 -4.800 2798.690 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.730 -4.800 894.290 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.290 -4.800 910.850 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.850 -4.800 927.410 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.410 -4.800 943.970 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.530 -4.800 977.090 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.090 -4.800 993.650 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.650 -4.800 1010.210 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.570 -4.800 712.130 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.210 -4.800 1026.770 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.330 -4.800 1059.890 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.890 -4.800 1076.450 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.450 -4.800 1093.010 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.010 -4.800 1109.570 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.130 -4.800 1142.690 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.690 -4.800 1159.250 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.250 -4.800 1175.810 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.930 -4.800 1225.490 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.490 -4.800 1242.050 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.050 -4.800 1258.610 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.610 -4.800 1275.170 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.730 -4.800 1308.290 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1324.290 -4.800 1324.850 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.850 -4.800 1341.410 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.690 -4.800 745.250 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1357.410 -4.800 1357.970 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1390.530 -4.800 1391.090 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.090 -4.800 1407.650 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1440.210 -4.800 1440.770 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.330 -4.800 1473.890 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.890 -4.800 1490.450 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.450 -4.800 1507.010 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.250 -4.800 761.810 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.010 -4.800 1523.570 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1556.130 -4.800 1556.690 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.250 -4.800 1589.810 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.810 -4.800 1606.370 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.370 -4.800 1622.930 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1638.930 -4.800 1639.490 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1655.490 -4.800 1656.050 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.050 -4.800 1672.610 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.810 -4.800 778.370 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1688.610 -4.800 1689.170 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1705.170 -4.800 1705.730 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.730 -4.800 1722.290 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.290 -4.800 1738.850 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.850 -4.800 1755.410 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.410 -4.800 1771.970 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.970 -4.800 1788.530 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1821.090 -4.800 1821.650 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1837.650 -4.800 1838.210 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.210 -4.800 1854.770 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.770 -4.800 1871.330 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.330 -4.800 1887.890 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.890 -4.800 1904.450 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1920.450 -4.800 1921.010 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1937.010 -4.800 1937.570 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.570 -4.800 1954.130 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1970.130 -4.800 1970.690 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1986.690 -4.800 1987.250 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.250 -4.800 2003.810 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.930 -4.800 811.490 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.810 -4.800 2020.370 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2052.930 -4.800 2053.490 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2069.490 -4.800 2070.050 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2086.050 -4.800 2086.610 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2102.610 -4.800 2103.170 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2119.170 -4.800 2119.730 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2135.730 -4.800 2136.290 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2152.290 -4.800 2152.850 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2168.850 -4.800 2169.410 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.490 -4.800 828.050 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2185.410 -4.800 2185.970 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.970 -4.800 2202.530 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.530 -4.800 2219.090 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2235.090 -4.800 2235.650 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2251.650 -4.800 2252.210 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.770 -4.800 2285.330 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.330 -4.800 2301.890 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2317.890 -4.800 2318.450 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2334.450 -4.800 2335.010 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.050 -4.800 844.610 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2809.170 -4.800 2809.730 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2814.690 -4.800 2815.250 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2820.210 -4.800 2820.770 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 -38.270 12.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 258.970 -38.270 262.070 21.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.970 -38.270 512.070 21.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 758.970 -38.270 762.070 21.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1008.970 -38.270 1012.070 21.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1258.970 -38.270 1262.070 21.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1508.970 -38.270 1512.070 21.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 1758.970 -38.270 1762.070 21.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2008.970 -38.270 2012.070 20.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 -38.270 2262.070 21.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2508.970 -38.270 2512.070 21.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 2758.970 -38.270 2762.070 21.435 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 14.330 2963.250 17.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 194.330 20.940 197.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 374.330 20.940 377.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 554.330 20.940 557.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 734.330 20.940 737.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 914.330 20.940 917.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1094.330 20.940 1097.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1274.330 20.940 1277.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1454.330 20.940 1457.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1634.330 20.940 1637.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1814.330 20.940 1817.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1994.330 20.940 1997.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2174.330 20.940 2177.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2354.330 20.940 2357.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2534.330 20.940 2537.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2714.330 20.940 2717.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2894.330 20.940 2897.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3074.330 20.940 3077.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3254.330 2963.250 3257.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3434.330 2963.250 3437.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 194.330 2963.250 197.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 374.330 2963.250 377.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 554.330 2963.250 557.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 734.330 2963.250 737.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 914.330 2963.250 917.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1094.330 2963.250 1097.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1274.330 2963.250 1277.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1454.330 2963.250 1457.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1634.330 2963.250 1637.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1814.330 2963.250 1817.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1994.330 2963.250 1997.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2174.330 2963.250 2177.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2354.330 2963.250 2357.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2534.330 2963.250 2537.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2714.330 2963.250 2717.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2894.330 2963.250 2897.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 3074.330 2963.250 3077.430 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2796.170 -38.270 2799.270 3557.950 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 2833.370 -38.270 2836.470 194.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 2833.370 661.680 2836.470 844.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2833.370 1311.760 2836.470 1494.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 2833.370 1961.840 2836.470 2144.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2833.370 2611.920 2836.470 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 88.730 2963.250 91.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3328.730 2963.250 3331.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 808.730 2963.250 811.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1348.730 2963.250 1351.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2068.730 2963.250 2071.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2788.730 2963.250 2791.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2968.730 2963.250 2971.830 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 3148.730 2963.250 3151.830 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2870.570 -38.270 2873.670 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 125.930 2963.250 129.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3365.930 2963.250 3369.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 305.930 2963.250 309.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 485.930 2963.250 489.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 665.930 2963.250 669.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 845.930 2963.250 849.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1025.930 2963.250 1029.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1205.930 2963.250 1209.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1385.930 2963.250 1389.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1565.930 2963.250 1569.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1745.930 2963.250 1749.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1925.930 2963.250 1929.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2105.930 2963.250 2109.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2285.930 2963.250 2289.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2465.930 2963.250 2469.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2645.930 2963.250 2649.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2825.930 2963.250 2829.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 3005.930 2963.250 3009.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 3185.930 2963.250 3189.030 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2851.970 -38.270 2855.070 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 107.330 2963.250 110.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3347.330 2963.250 3350.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 287.330 2963.250 290.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 467.330 2963.250 470.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 647.330 2963.250 650.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 827.330 2963.250 830.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1007.330 2963.250 1010.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1187.330 2963.250 1190.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1367.330 2963.250 1370.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1547.330 2963.250 1550.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1727.330 2963.250 1730.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1907.330 2963.250 1910.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2087.330 2963.250 2090.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2267.330 2963.250 2270.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2447.330 2963.250 2450.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2627.330 2963.250 2630.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2807.330 2963.250 2810.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2987.330 2963.250 2990.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 3167.330 2963.250 3170.430 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2889.170 -38.270 2892.270 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 144.530 2963.250 147.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3384.530 2963.250 3387.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 324.530 2963.250 327.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 504.530 2963.250 507.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 684.530 2963.250 687.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 864.530 2963.250 867.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1044.530 2963.250 1047.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1224.530 2963.250 1227.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1404.530 2963.250 1407.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1584.530 2963.250 1587.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1764.530 2963.250 1767.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1944.530 2963.250 1947.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2124.530 2963.250 2127.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2304.530 2963.250 2307.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2484.530 2963.250 2487.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2664.530 2963.250 2667.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2844.530 2963.250 2847.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 3024.530 2963.250 3027.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 3204.530 2963.250 3207.630 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2777.570 -38.270 2780.670 3557.950 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2814.770 -38.270 2817.870 194.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 2814.770 661.680 2817.870 844.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2814.770 1311.760 2817.870 1494.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 2814.770 1961.840 2817.870 2144.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2814.770 2611.920 2817.870 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 70.130 2963.250 73.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3310.130 2963.250 3313.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3490.130 2963.250 3493.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 790.130 2963.250 793.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 1330.130 2963.250 1333.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2050.130 2963.250 2053.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2770.130 2963.250 2773.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 2950.130 2963.250 2953.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 2331.020 3130.130 2963.250 3133.230 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.850 -4.800 99.410 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.370 -4.800 104.930 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.890 -4.800 110.450 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.970 -4.800 132.530 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.650 -4.800 320.210 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.210 -4.800 336.770 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.770 -4.800 353.330 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.330 -4.800 369.890 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.890 -4.800 386.450 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.450 -4.800 403.010 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.570 -4.800 436.130 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.130 -4.800 452.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.690 -4.800 469.250 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.050 -4.800 154.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.250 -4.800 485.810 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.810 -4.800 502.370 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.370 -4.800 518.930 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.930 -4.800 535.490 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.490 -4.800 552.050 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.050 -4.800 568.610 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.610 -4.800 585.170 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.170 -4.800 601.730 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.730 -4.800 618.290 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.290 -4.800 634.850 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.130 -4.800 176.690 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.410 -4.800 667.970 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.210 -4.800 198.770 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.290 -4.800 220.850 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.850 -4.800 237.410 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.410 -4.800 253.970 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.530 -4.800 287.090 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.090 -4.800 303.650 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.490 -4.800 138.050 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.170 -4.800 325.730 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.730 -4.800 342.290 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.290 -4.800 358.850 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.410 -4.800 391.970 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.970 -4.800 408.530 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.090 -4.800 441.650 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.210 -4.800 474.770 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.570 -4.800 160.130 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.770 -4.800 491.330 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.330 -4.800 507.890 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.890 -4.800 524.450 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.010 -4.800 557.570 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.130 -4.800 590.690 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.690 -4.800 607.250 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.250 -4.800 623.810 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.810 -4.800 640.370 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.650 -4.800 182.210 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.370 -4.800 656.930 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.930 -4.800 673.490 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.730 -4.800 204.290 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.810 -4.800 226.370 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.370 -4.800 242.930 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.930 -4.800 259.490 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.490 -4.800 276.050 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.610 -4.800 309.170 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.010 -4.800 143.570 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.690 -4.800 331.250 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.810 -4.800 364.370 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.370 -4.800 380.930 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.930 -4.800 397.490 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.490 -4.800 414.050 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.050 -4.800 430.610 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.610 -4.800 447.170 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.170 -4.800 463.730 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.730 -4.800 480.290 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.090 -4.800 165.650 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.850 -4.800 513.410 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.410 -4.800 529.970 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.970 -4.800 546.530 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.530 -4.800 563.090 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.090 -4.800 579.650 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.650 -4.800 596.210 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.210 -4.800 612.770 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.770 -4.800 629.330 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.330 -4.800 645.890 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.170 -4.800 187.730 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.890 -4.800 662.450 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.450 -4.800 679.010 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.330 -4.800 231.890 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.890 -4.800 248.450 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.450 -4.800 265.010 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.010 -4.800 281.570 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.570 -4.800 298.130 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.130 -4.800 314.690 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.530 -4.800 149.090 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.610 -4.800 171.170 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.770 -4.800 215.330 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 25.520 30.795 2894.080 3488.085 ;
      LAYER met1 ;
        RECT 25.520 30.640 2894.080 3515.220 ;
      LAYER met2 ;
        RECT 6.530 3517.320 42.450 3518.050 ;
        RECT 43.570 3517.320 123.410 3518.050 ;
        RECT 124.530 3517.320 204.370 3518.050 ;
        RECT 205.490 3517.320 285.330 3518.050 ;
        RECT 286.450 3517.320 366.290 3518.050 ;
        RECT 367.410 3517.320 447.250 3518.050 ;
        RECT 448.370 3517.320 528.210 3518.050 ;
        RECT 529.330 3517.320 609.170 3518.050 ;
        RECT 610.290 3517.320 690.130 3518.050 ;
        RECT 691.250 3517.320 771.090 3518.050 ;
        RECT 772.210 3517.320 852.050 3518.050 ;
        RECT 853.170 3517.320 933.010 3518.050 ;
        RECT 934.130 3517.320 1013.970 3518.050 ;
        RECT 1015.090 3517.320 1094.930 3518.050 ;
        RECT 1096.050 3517.320 1175.890 3518.050 ;
        RECT 1177.010 3517.320 1256.850 3518.050 ;
        RECT 1257.970 3517.320 1337.810 3518.050 ;
        RECT 1338.930 3517.320 1418.770 3518.050 ;
        RECT 1419.890 3517.320 1499.730 3518.050 ;
        RECT 1500.850 3517.320 1580.690 3518.050 ;
        RECT 1581.810 3517.320 1661.650 3518.050 ;
        RECT 1662.770 3517.320 1742.610 3518.050 ;
        RECT 1743.730 3517.320 1823.570 3518.050 ;
        RECT 1824.690 3517.320 1904.530 3518.050 ;
        RECT 1905.650 3517.320 1985.490 3518.050 ;
        RECT 1986.610 3517.320 2066.450 3518.050 ;
        RECT 2067.570 3517.320 2147.410 3518.050 ;
        RECT 2148.530 3517.320 2228.370 3518.050 ;
        RECT 2229.490 3517.320 2309.330 3518.050 ;
        RECT 2310.450 3517.320 2390.290 3518.050 ;
        RECT 2391.410 3517.320 2471.250 3518.050 ;
        RECT 2472.370 3517.320 2552.210 3518.050 ;
        RECT 2553.330 3517.320 2633.170 3518.050 ;
        RECT 2634.290 3517.320 2714.130 3518.050 ;
        RECT 2715.250 3517.320 2795.090 3518.050 ;
        RECT 2796.210 3517.320 2876.050 3518.050 ;
        RECT 2877.170 3517.320 2912.170 3518.050 ;
        RECT 6.530 2.680 2912.170 3517.320 ;
        RECT 6.530 2.400 98.570 2.680 ;
        RECT 99.690 2.400 104.090 2.680 ;
        RECT 105.210 2.400 109.610 2.680 ;
        RECT 110.730 2.400 115.130 2.680 ;
        RECT 116.250 2.400 120.650 2.680 ;
        RECT 121.770 2.400 126.170 2.680 ;
        RECT 127.290 2.400 131.690 2.680 ;
        RECT 132.810 2.400 137.210 2.680 ;
        RECT 138.330 2.400 142.730 2.680 ;
        RECT 143.850 2.400 148.250 2.680 ;
        RECT 149.370 2.400 153.770 2.680 ;
        RECT 154.890 2.400 159.290 2.680 ;
        RECT 160.410 2.400 164.810 2.680 ;
        RECT 165.930 2.400 170.330 2.680 ;
        RECT 171.450 2.400 175.850 2.680 ;
        RECT 176.970 2.400 181.370 2.680 ;
        RECT 182.490 2.400 186.890 2.680 ;
        RECT 188.010 2.400 192.410 2.680 ;
        RECT 193.530 2.400 197.930 2.680 ;
        RECT 199.050 2.400 203.450 2.680 ;
        RECT 204.570 2.400 208.970 2.680 ;
        RECT 210.090 2.400 214.490 2.680 ;
        RECT 215.610 2.400 220.010 2.680 ;
        RECT 221.130 2.400 225.530 2.680 ;
        RECT 226.650 2.400 231.050 2.680 ;
        RECT 232.170 2.400 236.570 2.680 ;
        RECT 237.690 2.400 242.090 2.680 ;
        RECT 243.210 2.400 247.610 2.680 ;
        RECT 248.730 2.400 253.130 2.680 ;
        RECT 254.250 2.400 258.650 2.680 ;
        RECT 259.770 2.400 264.170 2.680 ;
        RECT 265.290 2.400 269.690 2.680 ;
        RECT 270.810 2.400 275.210 2.680 ;
        RECT 276.330 2.400 280.730 2.680 ;
        RECT 281.850 2.400 286.250 2.680 ;
        RECT 287.370 2.400 291.770 2.680 ;
        RECT 292.890 2.400 297.290 2.680 ;
        RECT 298.410 2.400 302.810 2.680 ;
        RECT 303.930 2.400 308.330 2.680 ;
        RECT 309.450 2.400 313.850 2.680 ;
        RECT 314.970 2.400 319.370 2.680 ;
        RECT 320.490 2.400 324.890 2.680 ;
        RECT 326.010 2.400 330.410 2.680 ;
        RECT 331.530 2.400 335.930 2.680 ;
        RECT 337.050 2.400 341.450 2.680 ;
        RECT 342.570 2.400 346.970 2.680 ;
        RECT 348.090 2.400 352.490 2.680 ;
        RECT 353.610 2.400 358.010 2.680 ;
        RECT 359.130 2.400 363.530 2.680 ;
        RECT 364.650 2.400 369.050 2.680 ;
        RECT 370.170 2.400 374.570 2.680 ;
        RECT 375.690 2.400 380.090 2.680 ;
        RECT 381.210 2.400 385.610 2.680 ;
        RECT 386.730 2.400 391.130 2.680 ;
        RECT 392.250 2.400 396.650 2.680 ;
        RECT 397.770 2.400 402.170 2.680 ;
        RECT 403.290 2.400 407.690 2.680 ;
        RECT 408.810 2.400 413.210 2.680 ;
        RECT 414.330 2.400 418.730 2.680 ;
        RECT 419.850 2.400 424.250 2.680 ;
        RECT 425.370 2.400 429.770 2.680 ;
        RECT 430.890 2.400 435.290 2.680 ;
        RECT 436.410 2.400 440.810 2.680 ;
        RECT 441.930 2.400 446.330 2.680 ;
        RECT 447.450 2.400 451.850 2.680 ;
        RECT 452.970 2.400 457.370 2.680 ;
        RECT 458.490 2.400 462.890 2.680 ;
        RECT 464.010 2.400 468.410 2.680 ;
        RECT 469.530 2.400 473.930 2.680 ;
        RECT 475.050 2.400 479.450 2.680 ;
        RECT 480.570 2.400 484.970 2.680 ;
        RECT 486.090 2.400 490.490 2.680 ;
        RECT 491.610 2.400 496.010 2.680 ;
        RECT 497.130 2.400 501.530 2.680 ;
        RECT 502.650 2.400 507.050 2.680 ;
        RECT 508.170 2.400 512.570 2.680 ;
        RECT 513.690 2.400 518.090 2.680 ;
        RECT 519.210 2.400 523.610 2.680 ;
        RECT 524.730 2.400 529.130 2.680 ;
        RECT 530.250 2.400 534.650 2.680 ;
        RECT 535.770 2.400 540.170 2.680 ;
        RECT 541.290 2.400 545.690 2.680 ;
        RECT 546.810 2.400 551.210 2.680 ;
        RECT 552.330 2.400 556.730 2.680 ;
        RECT 557.850 2.400 562.250 2.680 ;
        RECT 563.370 2.400 567.770 2.680 ;
        RECT 568.890 2.400 573.290 2.680 ;
        RECT 574.410 2.400 578.810 2.680 ;
        RECT 579.930 2.400 584.330 2.680 ;
        RECT 585.450 2.400 589.850 2.680 ;
        RECT 590.970 2.400 595.370 2.680 ;
        RECT 596.490 2.400 600.890 2.680 ;
        RECT 602.010 2.400 606.410 2.680 ;
        RECT 607.530 2.400 611.930 2.680 ;
        RECT 613.050 2.400 617.450 2.680 ;
        RECT 618.570 2.400 622.970 2.680 ;
        RECT 624.090 2.400 628.490 2.680 ;
        RECT 629.610 2.400 634.010 2.680 ;
        RECT 635.130 2.400 639.530 2.680 ;
        RECT 640.650 2.400 645.050 2.680 ;
        RECT 646.170 2.400 650.570 2.680 ;
        RECT 651.690 2.400 656.090 2.680 ;
        RECT 657.210 2.400 661.610 2.680 ;
        RECT 662.730 2.400 667.130 2.680 ;
        RECT 668.250 2.400 672.650 2.680 ;
        RECT 673.770 2.400 678.170 2.680 ;
        RECT 679.290 2.400 683.690 2.680 ;
        RECT 684.810 2.400 689.210 2.680 ;
        RECT 690.330 2.400 694.730 2.680 ;
        RECT 695.850 2.400 700.250 2.680 ;
        RECT 701.370 2.400 705.770 2.680 ;
        RECT 706.890 2.400 711.290 2.680 ;
        RECT 712.410 2.400 716.810 2.680 ;
        RECT 717.930 2.400 722.330 2.680 ;
        RECT 723.450 2.400 727.850 2.680 ;
        RECT 728.970 2.400 733.370 2.680 ;
        RECT 734.490 2.400 738.890 2.680 ;
        RECT 740.010 2.400 744.410 2.680 ;
        RECT 745.530 2.400 749.930 2.680 ;
        RECT 751.050 2.400 755.450 2.680 ;
        RECT 756.570 2.400 760.970 2.680 ;
        RECT 762.090 2.400 766.490 2.680 ;
        RECT 767.610 2.400 772.010 2.680 ;
        RECT 773.130 2.400 777.530 2.680 ;
        RECT 778.650 2.400 783.050 2.680 ;
        RECT 784.170 2.400 788.570 2.680 ;
        RECT 789.690 2.400 794.090 2.680 ;
        RECT 795.210 2.400 799.610 2.680 ;
        RECT 800.730 2.400 805.130 2.680 ;
        RECT 806.250 2.400 810.650 2.680 ;
        RECT 811.770 2.400 816.170 2.680 ;
        RECT 817.290 2.400 821.690 2.680 ;
        RECT 822.810 2.400 827.210 2.680 ;
        RECT 828.330 2.400 832.730 2.680 ;
        RECT 833.850 2.400 838.250 2.680 ;
        RECT 839.370 2.400 843.770 2.680 ;
        RECT 844.890 2.400 849.290 2.680 ;
        RECT 850.410 2.400 854.810 2.680 ;
        RECT 855.930 2.400 860.330 2.680 ;
        RECT 861.450 2.400 865.850 2.680 ;
        RECT 866.970 2.400 871.370 2.680 ;
        RECT 872.490 2.400 876.890 2.680 ;
        RECT 878.010 2.400 882.410 2.680 ;
        RECT 883.530 2.400 887.930 2.680 ;
        RECT 889.050 2.400 893.450 2.680 ;
        RECT 894.570 2.400 898.970 2.680 ;
        RECT 900.090 2.400 904.490 2.680 ;
        RECT 905.610 2.400 910.010 2.680 ;
        RECT 911.130 2.400 915.530 2.680 ;
        RECT 916.650 2.400 921.050 2.680 ;
        RECT 922.170 2.400 926.570 2.680 ;
        RECT 927.690 2.400 932.090 2.680 ;
        RECT 933.210 2.400 937.610 2.680 ;
        RECT 938.730 2.400 943.130 2.680 ;
        RECT 944.250 2.400 948.650 2.680 ;
        RECT 949.770 2.400 954.170 2.680 ;
        RECT 955.290 2.400 959.690 2.680 ;
        RECT 960.810 2.400 965.210 2.680 ;
        RECT 966.330 2.400 970.730 2.680 ;
        RECT 971.850 2.400 976.250 2.680 ;
        RECT 977.370 2.400 981.770 2.680 ;
        RECT 982.890 2.400 987.290 2.680 ;
        RECT 988.410 2.400 992.810 2.680 ;
        RECT 993.930 2.400 998.330 2.680 ;
        RECT 999.450 2.400 1003.850 2.680 ;
        RECT 1004.970 2.400 1009.370 2.680 ;
        RECT 1010.490 2.400 1014.890 2.680 ;
        RECT 1016.010 2.400 1020.410 2.680 ;
        RECT 1021.530 2.400 1025.930 2.680 ;
        RECT 1027.050 2.400 1031.450 2.680 ;
        RECT 1032.570 2.400 1036.970 2.680 ;
        RECT 1038.090 2.400 1042.490 2.680 ;
        RECT 1043.610 2.400 1048.010 2.680 ;
        RECT 1049.130 2.400 1053.530 2.680 ;
        RECT 1054.650 2.400 1059.050 2.680 ;
        RECT 1060.170 2.400 1064.570 2.680 ;
        RECT 1065.690 2.400 1070.090 2.680 ;
        RECT 1071.210 2.400 1075.610 2.680 ;
        RECT 1076.730 2.400 1081.130 2.680 ;
        RECT 1082.250 2.400 1086.650 2.680 ;
        RECT 1087.770 2.400 1092.170 2.680 ;
        RECT 1093.290 2.400 1097.690 2.680 ;
        RECT 1098.810 2.400 1103.210 2.680 ;
        RECT 1104.330 2.400 1108.730 2.680 ;
        RECT 1109.850 2.400 1114.250 2.680 ;
        RECT 1115.370 2.400 1119.770 2.680 ;
        RECT 1120.890 2.400 1125.290 2.680 ;
        RECT 1126.410 2.400 1130.810 2.680 ;
        RECT 1131.930 2.400 1136.330 2.680 ;
        RECT 1137.450 2.400 1141.850 2.680 ;
        RECT 1142.970 2.400 1147.370 2.680 ;
        RECT 1148.490 2.400 1152.890 2.680 ;
        RECT 1154.010 2.400 1158.410 2.680 ;
        RECT 1159.530 2.400 1163.930 2.680 ;
        RECT 1165.050 2.400 1169.450 2.680 ;
        RECT 1170.570 2.400 1174.970 2.680 ;
        RECT 1176.090 2.400 1180.490 2.680 ;
        RECT 1181.610 2.400 1186.010 2.680 ;
        RECT 1187.130 2.400 1191.530 2.680 ;
        RECT 1192.650 2.400 1197.050 2.680 ;
        RECT 1198.170 2.400 1202.570 2.680 ;
        RECT 1203.690 2.400 1208.090 2.680 ;
        RECT 1209.210 2.400 1213.610 2.680 ;
        RECT 1214.730 2.400 1219.130 2.680 ;
        RECT 1220.250 2.400 1224.650 2.680 ;
        RECT 1225.770 2.400 1230.170 2.680 ;
        RECT 1231.290 2.400 1235.690 2.680 ;
        RECT 1236.810 2.400 1241.210 2.680 ;
        RECT 1242.330 2.400 1246.730 2.680 ;
        RECT 1247.850 2.400 1252.250 2.680 ;
        RECT 1253.370 2.400 1257.770 2.680 ;
        RECT 1258.890 2.400 1263.290 2.680 ;
        RECT 1264.410 2.400 1268.810 2.680 ;
        RECT 1269.930 2.400 1274.330 2.680 ;
        RECT 1275.450 2.400 1279.850 2.680 ;
        RECT 1280.970 2.400 1285.370 2.680 ;
        RECT 1286.490 2.400 1290.890 2.680 ;
        RECT 1292.010 2.400 1296.410 2.680 ;
        RECT 1297.530 2.400 1301.930 2.680 ;
        RECT 1303.050 2.400 1307.450 2.680 ;
        RECT 1308.570 2.400 1312.970 2.680 ;
        RECT 1314.090 2.400 1318.490 2.680 ;
        RECT 1319.610 2.400 1324.010 2.680 ;
        RECT 1325.130 2.400 1329.530 2.680 ;
        RECT 1330.650 2.400 1335.050 2.680 ;
        RECT 1336.170 2.400 1340.570 2.680 ;
        RECT 1341.690 2.400 1346.090 2.680 ;
        RECT 1347.210 2.400 1351.610 2.680 ;
        RECT 1352.730 2.400 1357.130 2.680 ;
        RECT 1358.250 2.400 1362.650 2.680 ;
        RECT 1363.770 2.400 1368.170 2.680 ;
        RECT 1369.290 2.400 1373.690 2.680 ;
        RECT 1374.810 2.400 1379.210 2.680 ;
        RECT 1380.330 2.400 1384.730 2.680 ;
        RECT 1385.850 2.400 1390.250 2.680 ;
        RECT 1391.370 2.400 1395.770 2.680 ;
        RECT 1396.890 2.400 1401.290 2.680 ;
        RECT 1402.410 2.400 1406.810 2.680 ;
        RECT 1407.930 2.400 1412.330 2.680 ;
        RECT 1413.450 2.400 1417.850 2.680 ;
        RECT 1418.970 2.400 1423.370 2.680 ;
        RECT 1424.490 2.400 1428.890 2.680 ;
        RECT 1430.010 2.400 1434.410 2.680 ;
        RECT 1435.530 2.400 1439.930 2.680 ;
        RECT 1441.050 2.400 1445.450 2.680 ;
        RECT 1446.570 2.400 1450.970 2.680 ;
        RECT 1452.090 2.400 1456.490 2.680 ;
        RECT 1457.610 2.400 1462.010 2.680 ;
        RECT 1463.130 2.400 1467.530 2.680 ;
        RECT 1468.650 2.400 1473.050 2.680 ;
        RECT 1474.170 2.400 1478.570 2.680 ;
        RECT 1479.690 2.400 1484.090 2.680 ;
        RECT 1485.210 2.400 1489.610 2.680 ;
        RECT 1490.730 2.400 1495.130 2.680 ;
        RECT 1496.250 2.400 1500.650 2.680 ;
        RECT 1501.770 2.400 1506.170 2.680 ;
        RECT 1507.290 2.400 1511.690 2.680 ;
        RECT 1512.810 2.400 1517.210 2.680 ;
        RECT 1518.330 2.400 1522.730 2.680 ;
        RECT 1523.850 2.400 1528.250 2.680 ;
        RECT 1529.370 2.400 1533.770 2.680 ;
        RECT 1534.890 2.400 1539.290 2.680 ;
        RECT 1540.410 2.400 1544.810 2.680 ;
        RECT 1545.930 2.400 1550.330 2.680 ;
        RECT 1551.450 2.400 1555.850 2.680 ;
        RECT 1556.970 2.400 1561.370 2.680 ;
        RECT 1562.490 2.400 1566.890 2.680 ;
        RECT 1568.010 2.400 1572.410 2.680 ;
        RECT 1573.530 2.400 1577.930 2.680 ;
        RECT 1579.050 2.400 1583.450 2.680 ;
        RECT 1584.570 2.400 1588.970 2.680 ;
        RECT 1590.090 2.400 1594.490 2.680 ;
        RECT 1595.610 2.400 1600.010 2.680 ;
        RECT 1601.130 2.400 1605.530 2.680 ;
        RECT 1606.650 2.400 1611.050 2.680 ;
        RECT 1612.170 2.400 1616.570 2.680 ;
        RECT 1617.690 2.400 1622.090 2.680 ;
        RECT 1623.210 2.400 1627.610 2.680 ;
        RECT 1628.730 2.400 1633.130 2.680 ;
        RECT 1634.250 2.400 1638.650 2.680 ;
        RECT 1639.770 2.400 1644.170 2.680 ;
        RECT 1645.290 2.400 1649.690 2.680 ;
        RECT 1650.810 2.400 1655.210 2.680 ;
        RECT 1656.330 2.400 1660.730 2.680 ;
        RECT 1661.850 2.400 1666.250 2.680 ;
        RECT 1667.370 2.400 1671.770 2.680 ;
        RECT 1672.890 2.400 1677.290 2.680 ;
        RECT 1678.410 2.400 1682.810 2.680 ;
        RECT 1683.930 2.400 1688.330 2.680 ;
        RECT 1689.450 2.400 1693.850 2.680 ;
        RECT 1694.970 2.400 1699.370 2.680 ;
        RECT 1700.490 2.400 1704.890 2.680 ;
        RECT 1706.010 2.400 1710.410 2.680 ;
        RECT 1711.530 2.400 1715.930 2.680 ;
        RECT 1717.050 2.400 1721.450 2.680 ;
        RECT 1722.570 2.400 1726.970 2.680 ;
        RECT 1728.090 2.400 1732.490 2.680 ;
        RECT 1733.610 2.400 1738.010 2.680 ;
        RECT 1739.130 2.400 1743.530 2.680 ;
        RECT 1744.650 2.400 1749.050 2.680 ;
        RECT 1750.170 2.400 1754.570 2.680 ;
        RECT 1755.690 2.400 1760.090 2.680 ;
        RECT 1761.210 2.400 1765.610 2.680 ;
        RECT 1766.730 2.400 1771.130 2.680 ;
        RECT 1772.250 2.400 1776.650 2.680 ;
        RECT 1777.770 2.400 1782.170 2.680 ;
        RECT 1783.290 2.400 1787.690 2.680 ;
        RECT 1788.810 2.400 1793.210 2.680 ;
        RECT 1794.330 2.400 1798.730 2.680 ;
        RECT 1799.850 2.400 1804.250 2.680 ;
        RECT 1805.370 2.400 1809.770 2.680 ;
        RECT 1810.890 2.400 1815.290 2.680 ;
        RECT 1816.410 2.400 1820.810 2.680 ;
        RECT 1821.930 2.400 1826.330 2.680 ;
        RECT 1827.450 2.400 1831.850 2.680 ;
        RECT 1832.970 2.400 1837.370 2.680 ;
        RECT 1838.490 2.400 1842.890 2.680 ;
        RECT 1844.010 2.400 1848.410 2.680 ;
        RECT 1849.530 2.400 1853.930 2.680 ;
        RECT 1855.050 2.400 1859.450 2.680 ;
        RECT 1860.570 2.400 1864.970 2.680 ;
        RECT 1866.090 2.400 1870.490 2.680 ;
        RECT 1871.610 2.400 1876.010 2.680 ;
        RECT 1877.130 2.400 1881.530 2.680 ;
        RECT 1882.650 2.400 1887.050 2.680 ;
        RECT 1888.170 2.400 1892.570 2.680 ;
        RECT 1893.690 2.400 1898.090 2.680 ;
        RECT 1899.210 2.400 1903.610 2.680 ;
        RECT 1904.730 2.400 1909.130 2.680 ;
        RECT 1910.250 2.400 1914.650 2.680 ;
        RECT 1915.770 2.400 1920.170 2.680 ;
        RECT 1921.290 2.400 1925.690 2.680 ;
        RECT 1926.810 2.400 1931.210 2.680 ;
        RECT 1932.330 2.400 1936.730 2.680 ;
        RECT 1937.850 2.400 1942.250 2.680 ;
        RECT 1943.370 2.400 1947.770 2.680 ;
        RECT 1948.890 2.400 1953.290 2.680 ;
        RECT 1954.410 2.400 1958.810 2.680 ;
        RECT 1959.930 2.400 1964.330 2.680 ;
        RECT 1965.450 2.400 1969.850 2.680 ;
        RECT 1970.970 2.400 1975.370 2.680 ;
        RECT 1976.490 2.400 1980.890 2.680 ;
        RECT 1982.010 2.400 1986.410 2.680 ;
        RECT 1987.530 2.400 1991.930 2.680 ;
        RECT 1993.050 2.400 1997.450 2.680 ;
        RECT 1998.570 2.400 2002.970 2.680 ;
        RECT 2004.090 2.400 2008.490 2.680 ;
        RECT 2009.610 2.400 2014.010 2.680 ;
        RECT 2015.130 2.400 2019.530 2.680 ;
        RECT 2020.650 2.400 2025.050 2.680 ;
        RECT 2026.170 2.400 2030.570 2.680 ;
        RECT 2031.690 2.400 2036.090 2.680 ;
        RECT 2037.210 2.400 2041.610 2.680 ;
        RECT 2042.730 2.400 2047.130 2.680 ;
        RECT 2048.250 2.400 2052.650 2.680 ;
        RECT 2053.770 2.400 2058.170 2.680 ;
        RECT 2059.290 2.400 2063.690 2.680 ;
        RECT 2064.810 2.400 2069.210 2.680 ;
        RECT 2070.330 2.400 2074.730 2.680 ;
        RECT 2075.850 2.400 2080.250 2.680 ;
        RECT 2081.370 2.400 2085.770 2.680 ;
        RECT 2086.890 2.400 2091.290 2.680 ;
        RECT 2092.410 2.400 2096.810 2.680 ;
        RECT 2097.930 2.400 2102.330 2.680 ;
        RECT 2103.450 2.400 2107.850 2.680 ;
        RECT 2108.970 2.400 2113.370 2.680 ;
        RECT 2114.490 2.400 2118.890 2.680 ;
        RECT 2120.010 2.400 2124.410 2.680 ;
        RECT 2125.530 2.400 2129.930 2.680 ;
        RECT 2131.050 2.400 2135.450 2.680 ;
        RECT 2136.570 2.400 2140.970 2.680 ;
        RECT 2142.090 2.400 2146.490 2.680 ;
        RECT 2147.610 2.400 2152.010 2.680 ;
        RECT 2153.130 2.400 2157.530 2.680 ;
        RECT 2158.650 2.400 2163.050 2.680 ;
        RECT 2164.170 2.400 2168.570 2.680 ;
        RECT 2169.690 2.400 2174.090 2.680 ;
        RECT 2175.210 2.400 2179.610 2.680 ;
        RECT 2180.730 2.400 2185.130 2.680 ;
        RECT 2186.250 2.400 2190.650 2.680 ;
        RECT 2191.770 2.400 2196.170 2.680 ;
        RECT 2197.290 2.400 2201.690 2.680 ;
        RECT 2202.810 2.400 2207.210 2.680 ;
        RECT 2208.330 2.400 2212.730 2.680 ;
        RECT 2213.850 2.400 2218.250 2.680 ;
        RECT 2219.370 2.400 2223.770 2.680 ;
        RECT 2224.890 2.400 2229.290 2.680 ;
        RECT 2230.410 2.400 2234.810 2.680 ;
        RECT 2235.930 2.400 2240.330 2.680 ;
        RECT 2241.450 2.400 2245.850 2.680 ;
        RECT 2246.970 2.400 2251.370 2.680 ;
        RECT 2252.490 2.400 2256.890 2.680 ;
        RECT 2258.010 2.400 2262.410 2.680 ;
        RECT 2263.530 2.400 2267.930 2.680 ;
        RECT 2269.050 2.400 2273.450 2.680 ;
        RECT 2274.570 2.400 2278.970 2.680 ;
        RECT 2280.090 2.400 2284.490 2.680 ;
        RECT 2285.610 2.400 2290.010 2.680 ;
        RECT 2291.130 2.400 2295.530 2.680 ;
        RECT 2296.650 2.400 2301.050 2.680 ;
        RECT 2302.170 2.400 2306.570 2.680 ;
        RECT 2307.690 2.400 2312.090 2.680 ;
        RECT 2313.210 2.400 2317.610 2.680 ;
        RECT 2318.730 2.400 2323.130 2.680 ;
        RECT 2324.250 2.400 2328.650 2.680 ;
        RECT 2329.770 2.400 2334.170 2.680 ;
        RECT 2335.290 2.400 2339.690 2.680 ;
        RECT 2340.810 2.400 2345.210 2.680 ;
        RECT 2346.330 2.400 2350.730 2.680 ;
        RECT 2351.850 2.400 2356.250 2.680 ;
        RECT 2357.370 2.400 2361.770 2.680 ;
        RECT 2362.890 2.400 2367.290 2.680 ;
        RECT 2368.410 2.400 2372.810 2.680 ;
        RECT 2373.930 2.400 2378.330 2.680 ;
        RECT 2379.450 2.400 2383.850 2.680 ;
        RECT 2384.970 2.400 2389.370 2.680 ;
        RECT 2390.490 2.400 2394.890 2.680 ;
        RECT 2396.010 2.400 2400.410 2.680 ;
        RECT 2401.530 2.400 2405.930 2.680 ;
        RECT 2407.050 2.400 2411.450 2.680 ;
        RECT 2412.570 2.400 2416.970 2.680 ;
        RECT 2418.090 2.400 2422.490 2.680 ;
        RECT 2423.610 2.400 2428.010 2.680 ;
        RECT 2429.130 2.400 2433.530 2.680 ;
        RECT 2434.650 2.400 2439.050 2.680 ;
        RECT 2440.170 2.400 2444.570 2.680 ;
        RECT 2445.690 2.400 2450.090 2.680 ;
        RECT 2451.210 2.400 2455.610 2.680 ;
        RECT 2456.730 2.400 2461.130 2.680 ;
        RECT 2462.250 2.400 2466.650 2.680 ;
        RECT 2467.770 2.400 2472.170 2.680 ;
        RECT 2473.290 2.400 2477.690 2.680 ;
        RECT 2478.810 2.400 2483.210 2.680 ;
        RECT 2484.330 2.400 2488.730 2.680 ;
        RECT 2489.850 2.400 2494.250 2.680 ;
        RECT 2495.370 2.400 2499.770 2.680 ;
        RECT 2500.890 2.400 2505.290 2.680 ;
        RECT 2506.410 2.400 2510.810 2.680 ;
        RECT 2511.930 2.400 2516.330 2.680 ;
        RECT 2517.450 2.400 2521.850 2.680 ;
        RECT 2522.970 2.400 2527.370 2.680 ;
        RECT 2528.490 2.400 2532.890 2.680 ;
        RECT 2534.010 2.400 2538.410 2.680 ;
        RECT 2539.530 2.400 2543.930 2.680 ;
        RECT 2545.050 2.400 2549.450 2.680 ;
        RECT 2550.570 2.400 2554.970 2.680 ;
        RECT 2556.090 2.400 2560.490 2.680 ;
        RECT 2561.610 2.400 2566.010 2.680 ;
        RECT 2567.130 2.400 2571.530 2.680 ;
        RECT 2572.650 2.400 2577.050 2.680 ;
        RECT 2578.170 2.400 2582.570 2.680 ;
        RECT 2583.690 2.400 2588.090 2.680 ;
        RECT 2589.210 2.400 2593.610 2.680 ;
        RECT 2594.730 2.400 2599.130 2.680 ;
        RECT 2600.250 2.400 2604.650 2.680 ;
        RECT 2605.770 2.400 2610.170 2.680 ;
        RECT 2611.290 2.400 2615.690 2.680 ;
        RECT 2616.810 2.400 2621.210 2.680 ;
        RECT 2622.330 2.400 2626.730 2.680 ;
        RECT 2627.850 2.400 2632.250 2.680 ;
        RECT 2633.370 2.400 2637.770 2.680 ;
        RECT 2638.890 2.400 2643.290 2.680 ;
        RECT 2644.410 2.400 2648.810 2.680 ;
        RECT 2649.930 2.400 2654.330 2.680 ;
        RECT 2655.450 2.400 2659.850 2.680 ;
        RECT 2660.970 2.400 2665.370 2.680 ;
        RECT 2666.490 2.400 2670.890 2.680 ;
        RECT 2672.010 2.400 2676.410 2.680 ;
        RECT 2677.530 2.400 2681.930 2.680 ;
        RECT 2683.050 2.400 2687.450 2.680 ;
        RECT 2688.570 2.400 2692.970 2.680 ;
        RECT 2694.090 2.400 2698.490 2.680 ;
        RECT 2699.610 2.400 2704.010 2.680 ;
        RECT 2705.130 2.400 2709.530 2.680 ;
        RECT 2710.650 2.400 2715.050 2.680 ;
        RECT 2716.170 2.400 2720.570 2.680 ;
        RECT 2721.690 2.400 2726.090 2.680 ;
        RECT 2727.210 2.400 2731.610 2.680 ;
        RECT 2732.730 2.400 2737.130 2.680 ;
        RECT 2738.250 2.400 2742.650 2.680 ;
        RECT 2743.770 2.400 2748.170 2.680 ;
        RECT 2749.290 2.400 2753.690 2.680 ;
        RECT 2754.810 2.400 2759.210 2.680 ;
        RECT 2760.330 2.400 2764.730 2.680 ;
        RECT 2765.850 2.400 2770.250 2.680 ;
        RECT 2771.370 2.400 2775.770 2.680 ;
        RECT 2776.890 2.400 2781.290 2.680 ;
        RECT 2782.410 2.400 2786.810 2.680 ;
        RECT 2787.930 2.400 2792.330 2.680 ;
        RECT 2793.450 2.400 2797.850 2.680 ;
        RECT 2798.970 2.400 2803.370 2.680 ;
        RECT 2804.490 2.400 2808.890 2.680 ;
        RECT 2810.010 2.400 2814.410 2.680 ;
        RECT 2815.530 2.400 2819.930 2.680 ;
        RECT 2821.050 2.400 2912.170 2.680 ;
      LAYER met3 ;
        RECT 1.230 3475.460 2917.930 3488.165 ;
        RECT 1.230 3473.460 2917.200 3475.460 ;
        RECT 1.230 3472.740 2917.930 3473.460 ;
        RECT 2.800 3470.740 2917.930 3472.740 ;
        RECT 1.230 3409.500 2917.930 3470.740 ;
        RECT 1.230 3408.140 2917.200 3409.500 ;
        RECT 2.800 3407.500 2917.200 3408.140 ;
        RECT 2.800 3406.140 2917.930 3407.500 ;
        RECT 1.230 3343.540 2917.930 3406.140 ;
        RECT 2.800 3341.540 2917.200 3343.540 ;
        RECT 1.230 3278.940 2917.930 3341.540 ;
        RECT 2.800 3277.580 2917.930 3278.940 ;
        RECT 2.800 3276.940 2917.200 3277.580 ;
        RECT 1.230 3275.580 2917.200 3276.940 ;
        RECT 1.230 3214.340 2917.930 3275.580 ;
        RECT 2.800 3212.340 2917.930 3214.340 ;
        RECT 1.230 3211.620 2917.930 3212.340 ;
        RECT 1.230 3209.620 2917.200 3211.620 ;
        RECT 1.230 3149.740 2917.930 3209.620 ;
        RECT 2.800 3147.740 2917.930 3149.740 ;
        RECT 1.230 3145.660 2917.930 3147.740 ;
        RECT 1.230 3143.660 2917.200 3145.660 ;
        RECT 1.230 3085.140 2917.930 3143.660 ;
        RECT 2.800 3083.140 2917.930 3085.140 ;
        RECT 1.230 3079.700 2917.930 3083.140 ;
        RECT 1.230 3077.700 2917.200 3079.700 ;
        RECT 1.230 3020.540 2917.930 3077.700 ;
        RECT 2.800 3018.540 2917.930 3020.540 ;
        RECT 1.230 3013.740 2917.930 3018.540 ;
        RECT 1.230 3011.740 2917.200 3013.740 ;
        RECT 1.230 2955.940 2917.930 3011.740 ;
        RECT 2.800 2953.940 2917.930 2955.940 ;
        RECT 1.230 2947.780 2917.930 2953.940 ;
        RECT 1.230 2945.780 2917.200 2947.780 ;
        RECT 1.230 2891.340 2917.930 2945.780 ;
        RECT 2.800 2889.340 2917.930 2891.340 ;
        RECT 1.230 2881.820 2917.930 2889.340 ;
        RECT 1.230 2879.820 2917.200 2881.820 ;
        RECT 1.230 2826.740 2917.930 2879.820 ;
        RECT 2.800 2824.740 2917.930 2826.740 ;
        RECT 1.230 2815.860 2917.930 2824.740 ;
        RECT 1.230 2813.860 2917.200 2815.860 ;
        RECT 1.230 2762.140 2917.930 2813.860 ;
        RECT 2.800 2760.140 2917.930 2762.140 ;
        RECT 1.230 2749.900 2917.930 2760.140 ;
        RECT 1.230 2747.900 2917.200 2749.900 ;
        RECT 1.230 2697.540 2917.930 2747.900 ;
        RECT 2.800 2695.540 2917.930 2697.540 ;
        RECT 1.230 2683.940 2917.930 2695.540 ;
        RECT 1.230 2681.940 2917.200 2683.940 ;
        RECT 1.230 2632.940 2917.930 2681.940 ;
        RECT 2.800 2630.940 2917.930 2632.940 ;
        RECT 1.230 2617.980 2917.930 2630.940 ;
        RECT 1.230 2615.980 2917.200 2617.980 ;
        RECT 1.230 2568.340 2917.930 2615.980 ;
        RECT 2.800 2566.340 2917.930 2568.340 ;
        RECT 1.230 2552.020 2917.930 2566.340 ;
        RECT 1.230 2550.020 2917.200 2552.020 ;
        RECT 1.230 2503.740 2917.930 2550.020 ;
        RECT 2.800 2501.740 2917.930 2503.740 ;
        RECT 1.230 2486.060 2917.930 2501.740 ;
        RECT 1.230 2484.060 2917.200 2486.060 ;
        RECT 1.230 2439.140 2917.930 2484.060 ;
        RECT 2.800 2437.140 2917.930 2439.140 ;
        RECT 1.230 2420.100 2917.930 2437.140 ;
        RECT 1.230 2418.100 2917.200 2420.100 ;
        RECT 1.230 2374.540 2917.930 2418.100 ;
        RECT 2.800 2372.540 2917.930 2374.540 ;
        RECT 1.230 2354.140 2917.930 2372.540 ;
        RECT 1.230 2352.140 2917.200 2354.140 ;
        RECT 1.230 2309.940 2917.930 2352.140 ;
        RECT 2.800 2307.940 2917.930 2309.940 ;
        RECT 1.230 2288.180 2917.930 2307.940 ;
        RECT 1.230 2286.180 2917.200 2288.180 ;
        RECT 1.230 2245.340 2917.930 2286.180 ;
        RECT 2.800 2243.340 2917.930 2245.340 ;
        RECT 1.230 2222.220 2917.930 2243.340 ;
        RECT 1.230 2220.220 2917.200 2222.220 ;
        RECT 1.230 2180.740 2917.930 2220.220 ;
        RECT 2.800 2178.740 2917.930 2180.740 ;
        RECT 1.230 2156.260 2917.930 2178.740 ;
        RECT 1.230 2154.260 2917.200 2156.260 ;
        RECT 1.230 2116.140 2917.930 2154.260 ;
        RECT 2.800 2114.140 2917.930 2116.140 ;
        RECT 1.230 2090.300 2917.930 2114.140 ;
        RECT 1.230 2088.300 2917.200 2090.300 ;
        RECT 1.230 2051.540 2917.930 2088.300 ;
        RECT 2.800 2049.540 2917.930 2051.540 ;
        RECT 1.230 2024.340 2917.930 2049.540 ;
        RECT 1.230 2022.340 2917.200 2024.340 ;
        RECT 1.230 1986.940 2917.930 2022.340 ;
        RECT 2.800 1984.940 2917.930 1986.940 ;
        RECT 1.230 1958.380 2917.930 1984.940 ;
        RECT 1.230 1956.380 2917.200 1958.380 ;
        RECT 1.230 1922.340 2917.930 1956.380 ;
        RECT 2.800 1920.340 2917.930 1922.340 ;
        RECT 1.230 1892.420 2917.930 1920.340 ;
        RECT 1.230 1890.420 2917.200 1892.420 ;
        RECT 1.230 1857.740 2917.930 1890.420 ;
        RECT 2.800 1855.740 2917.930 1857.740 ;
        RECT 1.230 1826.460 2917.930 1855.740 ;
        RECT 1.230 1824.460 2917.200 1826.460 ;
        RECT 1.230 1793.140 2917.930 1824.460 ;
        RECT 2.800 1791.140 2917.930 1793.140 ;
        RECT 1.230 1760.500 2917.930 1791.140 ;
        RECT 1.230 1758.500 2917.200 1760.500 ;
        RECT 1.230 1728.540 2917.930 1758.500 ;
        RECT 2.800 1726.540 2917.930 1728.540 ;
        RECT 1.230 1694.540 2917.930 1726.540 ;
        RECT 1.230 1692.540 2917.200 1694.540 ;
        RECT 1.230 1663.940 2917.930 1692.540 ;
        RECT 2.800 1661.940 2917.930 1663.940 ;
        RECT 1.230 1628.580 2917.930 1661.940 ;
        RECT 1.230 1626.580 2917.200 1628.580 ;
        RECT 1.230 1599.340 2917.930 1626.580 ;
        RECT 2.800 1597.340 2917.930 1599.340 ;
        RECT 1.230 1562.620 2917.930 1597.340 ;
        RECT 1.230 1560.620 2917.200 1562.620 ;
        RECT 1.230 1534.740 2917.930 1560.620 ;
        RECT 2.800 1532.740 2917.930 1534.740 ;
        RECT 1.230 1496.660 2917.930 1532.740 ;
        RECT 1.230 1494.660 2917.200 1496.660 ;
        RECT 1.230 1470.140 2917.930 1494.660 ;
        RECT 2.800 1468.140 2917.930 1470.140 ;
        RECT 1.230 1430.700 2917.930 1468.140 ;
        RECT 1.230 1428.700 2917.200 1430.700 ;
        RECT 1.230 1405.540 2917.930 1428.700 ;
        RECT 2.800 1403.540 2917.930 1405.540 ;
        RECT 1.230 1364.740 2917.930 1403.540 ;
        RECT 1.230 1362.740 2917.200 1364.740 ;
        RECT 1.230 1340.940 2917.930 1362.740 ;
        RECT 2.800 1338.940 2917.930 1340.940 ;
        RECT 1.230 1298.780 2917.930 1338.940 ;
        RECT 1.230 1296.780 2917.200 1298.780 ;
        RECT 1.230 1276.340 2917.930 1296.780 ;
        RECT 2.800 1274.340 2917.930 1276.340 ;
        RECT 1.230 1232.820 2917.930 1274.340 ;
        RECT 1.230 1230.820 2917.200 1232.820 ;
        RECT 1.230 1211.740 2917.930 1230.820 ;
        RECT 2.800 1209.740 2917.930 1211.740 ;
        RECT 1.230 1166.860 2917.930 1209.740 ;
        RECT 1.230 1164.860 2917.200 1166.860 ;
        RECT 1.230 1147.140 2917.930 1164.860 ;
        RECT 2.800 1145.140 2917.930 1147.140 ;
        RECT 1.230 1100.900 2917.930 1145.140 ;
        RECT 1.230 1098.900 2917.200 1100.900 ;
        RECT 1.230 1082.540 2917.930 1098.900 ;
        RECT 2.800 1080.540 2917.930 1082.540 ;
        RECT 1.230 1034.940 2917.930 1080.540 ;
        RECT 1.230 1032.940 2917.200 1034.940 ;
        RECT 1.230 1017.940 2917.930 1032.940 ;
        RECT 2.800 1015.940 2917.930 1017.940 ;
        RECT 1.230 968.980 2917.930 1015.940 ;
        RECT 1.230 966.980 2917.200 968.980 ;
        RECT 1.230 953.340 2917.930 966.980 ;
        RECT 2.800 951.340 2917.930 953.340 ;
        RECT 1.230 903.020 2917.930 951.340 ;
        RECT 1.230 901.020 2917.200 903.020 ;
        RECT 1.230 888.740 2917.930 901.020 ;
        RECT 2.800 886.740 2917.930 888.740 ;
        RECT 1.230 837.060 2917.930 886.740 ;
        RECT 1.230 835.060 2917.200 837.060 ;
        RECT 1.230 824.140 2917.930 835.060 ;
        RECT 2.800 822.140 2917.930 824.140 ;
        RECT 1.230 771.100 2917.930 822.140 ;
        RECT 1.230 769.100 2917.200 771.100 ;
        RECT 1.230 759.540 2917.930 769.100 ;
        RECT 2.800 757.540 2917.930 759.540 ;
        RECT 1.230 705.140 2917.930 757.540 ;
        RECT 1.230 703.140 2917.200 705.140 ;
        RECT 1.230 694.940 2917.930 703.140 ;
        RECT 2.800 692.940 2917.930 694.940 ;
        RECT 1.230 639.180 2917.930 692.940 ;
        RECT 1.230 637.180 2917.200 639.180 ;
        RECT 1.230 630.340 2917.930 637.180 ;
        RECT 2.800 628.340 2917.930 630.340 ;
        RECT 1.230 573.220 2917.930 628.340 ;
        RECT 1.230 571.220 2917.200 573.220 ;
        RECT 1.230 565.740 2917.930 571.220 ;
        RECT 2.800 563.740 2917.930 565.740 ;
        RECT 1.230 507.260 2917.930 563.740 ;
        RECT 1.230 505.260 2917.200 507.260 ;
        RECT 1.230 501.140 2917.930 505.260 ;
        RECT 2.800 499.140 2917.930 501.140 ;
        RECT 1.230 441.300 2917.930 499.140 ;
        RECT 1.230 439.300 2917.200 441.300 ;
        RECT 1.230 436.540 2917.930 439.300 ;
        RECT 2.800 434.540 2917.930 436.540 ;
        RECT 1.230 375.340 2917.930 434.540 ;
        RECT 1.230 373.340 2917.200 375.340 ;
        RECT 1.230 371.940 2917.930 373.340 ;
        RECT 2.800 369.940 2917.930 371.940 ;
        RECT 1.230 309.380 2917.930 369.940 ;
        RECT 1.230 307.380 2917.200 309.380 ;
        RECT 1.230 307.340 2917.930 307.380 ;
        RECT 2.800 305.340 2917.930 307.340 ;
        RECT 1.230 243.420 2917.930 305.340 ;
        RECT 1.230 242.740 2917.200 243.420 ;
        RECT 2.800 241.420 2917.200 242.740 ;
        RECT 2.800 240.740 2917.930 241.420 ;
        RECT 1.230 178.140 2917.930 240.740 ;
        RECT 2.800 177.460 2917.930 178.140 ;
        RECT 2.800 176.140 2917.200 177.460 ;
        RECT 1.230 175.460 2917.200 176.140 ;
        RECT 1.230 113.540 2917.930 175.460 ;
        RECT 2.800 111.540 2917.930 113.540 ;
        RECT 1.230 111.500 2917.930 111.540 ;
        RECT 1.230 109.500 2917.200 111.500 ;
        RECT 1.230 48.940 2917.930 109.500 ;
        RECT 2.800 46.940 2917.930 48.940 ;
        RECT 1.230 45.540 2917.930 46.940 ;
        RECT 1.230 43.540 2917.200 45.540 ;
        RECT 1.230 30.715 2917.930 43.540 ;
      LAYER met4 ;
        RECT 28.970 30.640 2777.170 3488.240 ;
        RECT 2781.070 30.640 2795.770 3488.240 ;
        RECT 2799.670 2611.520 2814.370 3488.240 ;
        RECT 2818.270 2611.520 2832.970 3488.240 ;
        RECT 2836.870 2611.520 2839.970 3488.240 ;
        RECT 2799.670 2144.960 2839.970 2611.520 ;
        RECT 2799.670 1961.440 2814.370 2144.960 ;
        RECT 2818.270 1961.440 2832.970 2144.960 ;
        RECT 2836.870 1961.440 2839.970 2144.960 ;
        RECT 2799.670 1494.880 2839.970 1961.440 ;
        RECT 2799.670 1311.360 2814.370 1494.880 ;
        RECT 2818.270 1311.360 2832.970 1494.880 ;
        RECT 2836.870 1311.360 2839.970 1494.880 ;
        RECT 2799.670 844.800 2839.970 1311.360 ;
        RECT 2799.670 661.280 2814.370 844.800 ;
        RECT 2818.270 661.280 2832.970 844.800 ;
        RECT 2836.870 661.280 2839.970 844.800 ;
        RECT 2799.670 194.720 2839.970 661.280 ;
        RECT 2799.670 30.640 2814.370 194.720 ;
        RECT 2818.270 30.640 2832.970 194.720 ;
        RECT 2836.870 30.640 2839.970 194.720 ;
      LAYER met5 ;
        RECT 25.280 3439.030 2894.320 3476.030 ;
        RECT 25.280 3389.230 2894.320 3432.730 ;
        RECT 25.280 3370.630 2894.320 3382.930 ;
        RECT 25.280 3352.030 2894.320 3364.330 ;
        RECT 25.280 3333.430 2894.320 3345.730 ;
        RECT 25.280 3314.830 2894.320 3327.130 ;
        RECT 25.280 3259.030 2894.320 3308.530 ;
        RECT 25.280 3209.230 2894.320 3252.730 ;
        RECT 25.280 3202.930 2329.420 3209.230 ;
        RECT 25.280 3190.630 2894.320 3202.930 ;
        RECT 25.280 3184.330 2329.420 3190.630 ;
        RECT 25.280 3172.030 2894.320 3184.330 ;
        RECT 25.280 3165.730 2329.420 3172.030 ;
        RECT 25.280 3153.430 2894.320 3165.730 ;
        RECT 25.280 3147.130 2329.420 3153.430 ;
        RECT 25.280 3134.830 2894.320 3147.130 ;
        RECT 25.280 3128.530 2329.420 3134.830 ;
        RECT 25.280 3079.030 2894.320 3128.530 ;
        RECT 25.280 3072.730 2329.420 3079.030 ;
        RECT 25.280 3029.230 2894.320 3072.730 ;
        RECT 25.280 3022.930 2329.420 3029.230 ;
        RECT 25.280 3010.630 2894.320 3022.930 ;
        RECT 25.280 3004.330 2329.420 3010.630 ;
        RECT 25.280 2992.030 2894.320 3004.330 ;
        RECT 25.280 2985.730 2329.420 2992.030 ;
        RECT 25.280 2973.430 2894.320 2985.730 ;
        RECT 25.280 2967.130 2329.420 2973.430 ;
        RECT 25.280 2954.830 2894.320 2967.130 ;
        RECT 25.280 2948.530 2329.420 2954.830 ;
        RECT 25.280 2899.030 2894.320 2948.530 ;
        RECT 25.280 2892.730 2329.420 2899.030 ;
        RECT 25.280 2849.230 2894.320 2892.730 ;
        RECT 25.280 2842.930 2329.420 2849.230 ;
        RECT 25.280 2830.630 2894.320 2842.930 ;
        RECT 25.280 2824.330 2329.420 2830.630 ;
        RECT 25.280 2812.030 2894.320 2824.330 ;
        RECT 25.280 2805.730 2329.420 2812.030 ;
        RECT 25.280 2793.430 2894.320 2805.730 ;
        RECT 25.280 2787.130 2329.420 2793.430 ;
        RECT 25.280 2774.830 2894.320 2787.130 ;
        RECT 25.280 2768.530 2329.420 2774.830 ;
        RECT 25.280 2719.030 2894.320 2768.530 ;
        RECT 25.280 2712.730 2329.420 2719.030 ;
        RECT 25.280 2669.230 2894.320 2712.730 ;
        RECT 25.280 2662.930 2329.420 2669.230 ;
        RECT 25.280 2650.630 2894.320 2662.930 ;
        RECT 25.280 2644.330 2329.420 2650.630 ;
        RECT 25.280 2632.030 2894.320 2644.330 ;
        RECT 25.280 2625.730 2329.420 2632.030 ;
        RECT 25.280 2539.030 2894.320 2625.730 ;
        RECT 25.280 2532.730 2329.420 2539.030 ;
        RECT 25.280 2489.230 2894.320 2532.730 ;
        RECT 25.280 2482.930 2329.420 2489.230 ;
        RECT 25.280 2470.630 2894.320 2482.930 ;
        RECT 25.280 2464.330 2329.420 2470.630 ;
        RECT 25.280 2452.030 2894.320 2464.330 ;
        RECT 25.280 2445.730 2329.420 2452.030 ;
        RECT 25.280 2359.030 2894.320 2445.730 ;
        RECT 25.280 2352.730 2329.420 2359.030 ;
        RECT 25.280 2309.230 2894.320 2352.730 ;
        RECT 25.280 2302.930 2329.420 2309.230 ;
        RECT 25.280 2290.630 2894.320 2302.930 ;
        RECT 25.280 2284.330 2329.420 2290.630 ;
        RECT 25.280 2272.030 2894.320 2284.330 ;
        RECT 25.280 2265.730 2329.420 2272.030 ;
        RECT 25.280 2179.030 2894.320 2265.730 ;
        RECT 25.280 2172.730 2329.420 2179.030 ;
        RECT 25.280 2129.230 2894.320 2172.730 ;
        RECT 25.280 2122.930 2329.420 2129.230 ;
        RECT 25.280 2110.630 2894.320 2122.930 ;
        RECT 25.280 2104.330 2329.420 2110.630 ;
        RECT 25.280 2092.030 2894.320 2104.330 ;
        RECT 25.280 2085.730 2329.420 2092.030 ;
        RECT 25.280 2073.430 2894.320 2085.730 ;
        RECT 25.280 2067.130 2329.420 2073.430 ;
        RECT 25.280 2054.830 2894.320 2067.130 ;
        RECT 25.280 2048.530 2329.420 2054.830 ;
        RECT 25.280 1999.030 2894.320 2048.530 ;
        RECT 25.280 1992.730 2329.420 1999.030 ;
        RECT 25.280 1949.230 2894.320 1992.730 ;
        RECT 25.280 1942.930 2329.420 1949.230 ;
        RECT 25.280 1930.630 2894.320 1942.930 ;
        RECT 25.280 1924.330 2329.420 1930.630 ;
        RECT 25.280 1912.030 2894.320 1924.330 ;
        RECT 25.280 1905.730 2329.420 1912.030 ;
        RECT 25.280 1819.030 2894.320 1905.730 ;
        RECT 25.280 1812.730 2329.420 1819.030 ;
        RECT 25.280 1769.230 2894.320 1812.730 ;
        RECT 25.280 1762.930 2329.420 1769.230 ;
        RECT 25.280 1750.630 2894.320 1762.930 ;
        RECT 25.280 1744.330 2329.420 1750.630 ;
        RECT 25.280 1732.030 2894.320 1744.330 ;
        RECT 25.280 1725.730 2329.420 1732.030 ;
        RECT 25.280 1639.030 2894.320 1725.730 ;
        RECT 25.280 1632.730 2329.420 1639.030 ;
        RECT 25.280 1589.230 2894.320 1632.730 ;
        RECT 25.280 1582.930 2329.420 1589.230 ;
        RECT 25.280 1570.630 2894.320 1582.930 ;
        RECT 25.280 1564.330 2329.420 1570.630 ;
        RECT 25.280 1552.030 2894.320 1564.330 ;
        RECT 25.280 1545.730 2329.420 1552.030 ;
        RECT 25.280 1459.030 2894.320 1545.730 ;
        RECT 25.280 1452.730 2329.420 1459.030 ;
        RECT 25.280 1409.230 2894.320 1452.730 ;
        RECT 25.280 1402.930 2329.420 1409.230 ;
        RECT 25.280 1390.630 2894.320 1402.930 ;
        RECT 25.280 1384.330 2329.420 1390.630 ;
        RECT 25.280 1372.030 2894.320 1384.330 ;
        RECT 25.280 1365.730 2329.420 1372.030 ;
        RECT 25.280 1353.430 2894.320 1365.730 ;
        RECT 25.280 1347.130 2329.420 1353.430 ;
        RECT 25.280 1334.830 2894.320 1347.130 ;
        RECT 25.280 1328.530 2329.420 1334.830 ;
        RECT 25.280 1279.030 2894.320 1328.530 ;
        RECT 25.280 1272.730 2329.420 1279.030 ;
        RECT 25.280 1229.230 2894.320 1272.730 ;
        RECT 25.280 1222.930 2329.420 1229.230 ;
        RECT 25.280 1210.630 2894.320 1222.930 ;
        RECT 25.280 1204.330 2329.420 1210.630 ;
        RECT 25.280 1192.030 2894.320 1204.330 ;
        RECT 25.280 1185.730 2329.420 1192.030 ;
        RECT 25.280 1099.030 2894.320 1185.730 ;
        RECT 25.280 1092.730 2329.420 1099.030 ;
        RECT 25.280 1049.230 2894.320 1092.730 ;
        RECT 25.280 1042.930 2329.420 1049.230 ;
        RECT 25.280 1030.630 2894.320 1042.930 ;
        RECT 25.280 1024.330 2329.420 1030.630 ;
        RECT 25.280 1012.030 2894.320 1024.330 ;
        RECT 25.280 1005.730 2329.420 1012.030 ;
        RECT 25.280 919.030 2894.320 1005.730 ;
        RECT 25.280 912.730 2329.420 919.030 ;
        RECT 25.280 869.230 2894.320 912.730 ;
        RECT 25.280 862.930 2329.420 869.230 ;
        RECT 25.280 850.630 2894.320 862.930 ;
        RECT 25.280 844.330 2329.420 850.630 ;
        RECT 25.280 832.030 2894.320 844.330 ;
        RECT 25.280 825.730 2329.420 832.030 ;
        RECT 25.280 813.430 2894.320 825.730 ;
        RECT 25.280 807.130 2329.420 813.430 ;
        RECT 25.280 794.830 2894.320 807.130 ;
        RECT 25.280 788.530 2329.420 794.830 ;
        RECT 25.280 739.030 2894.320 788.530 ;
        RECT 25.280 732.730 2329.420 739.030 ;
        RECT 25.280 689.230 2894.320 732.730 ;
        RECT 25.280 682.930 2329.420 689.230 ;
        RECT 25.280 670.630 2894.320 682.930 ;
        RECT 25.280 664.330 2329.420 670.630 ;
        RECT 25.280 652.030 2894.320 664.330 ;
        RECT 25.280 645.730 2329.420 652.030 ;
        RECT 25.280 559.030 2894.320 645.730 ;
        RECT 25.280 552.730 2329.420 559.030 ;
        RECT 25.280 509.230 2894.320 552.730 ;
        RECT 25.280 502.930 2329.420 509.230 ;
        RECT 25.280 490.630 2894.320 502.930 ;
        RECT 25.280 484.330 2329.420 490.630 ;
        RECT 25.280 472.030 2894.320 484.330 ;
        RECT 25.280 465.730 2329.420 472.030 ;
        RECT 25.280 379.030 2894.320 465.730 ;
        RECT 25.280 372.730 2329.420 379.030 ;
        RECT 25.280 329.230 2894.320 372.730 ;
        RECT 25.280 322.930 2329.420 329.230 ;
        RECT 25.280 310.630 2894.320 322.930 ;
        RECT 25.280 304.330 2329.420 310.630 ;
        RECT 25.280 292.030 2894.320 304.330 ;
        RECT 25.280 285.730 2329.420 292.030 ;
        RECT 25.280 199.030 2894.320 285.730 ;
        RECT 25.280 192.730 2329.420 199.030 ;
        RECT 25.280 149.230 2894.320 192.730 ;
        RECT 25.280 130.630 2894.320 142.930 ;
        RECT 25.280 112.030 2894.320 124.330 ;
        RECT 25.280 93.430 2894.320 105.730 ;
        RECT 25.280 74.830 2894.320 87.130 ;
        RECT 25.280 34.330 2894.320 68.530 ;
  END
END user_project_wrapper
END LIBRARY

